{ 16'sh_0001, 16'sh_0003, 16'sh_0005, 16'sh_000a, 16'sh_0014, 16'sh_0029, 16'sh_0051, 16'sh_00a3, 16'sh_0146, 16'sh_028c, 16'sh_0517, 16'sh_0a2c, 16'sh_1444, 16'sh_27ed, 16'sh_4b90, 16'sh_8000 }
