{ 9'sh_001, 9'sh_003, 9'sh_005, 9'sh_00a, 9'sh_014, 9'sh_029, 9'sh_050, 9'sh_097, 9'sh_100 }
