16'd237,
16'd257,
16'd276,
16'd296,
16'd316,
16'd336,
16'd356,
16'd375,
16'd395,
16'd415,
16'd478,
16'd502,
16'd526,
16'd550,
16'd574,
16'd597,
16'd621,
16'd645,
16'd669,
16'd692,
16'd716,
16'd740,
16'd764,
16'd787,
16'd811,
16'd835,
16'd859,
16'd883,
16'd906,
16'd930,
16'd954,
16'd978,
16'd1001,
16'd1025,
16'd1049,
16'd1073,
16'd1097,
16'd1120,
16'd1144,
16'd1168,
16'd1192,
16'd1215,
16'd1239,
16'd1263,
16'd1554,
16'd1584,
16'd1614,
16'd1643,
16'd1673,
16'd1703,
16'd1732,
16'd1762,
16'd1792,
16'd1822,
16'd1851,
16'd1881,
16'd1911,
16'd2515,
16'd2555,
16'd2594,
16'd2634,
16'd2674,
16'd3961,
16'd7825
