{ 24'sh_000001, 24'sh_000003, 24'sh_000005, 24'sh_00000a, 24'sh_000014, 24'sh_000029, 24'sh_000051, 24'sh_0000a3, 24'sh_000146, 24'sh_00028c, 24'sh_000518, 24'sh_000a30, 24'sh_00145f, 24'sh_0028be, 24'sh_00517d, 24'sh_00a2f9, 24'sh_0145f1, 24'sh_028bd8, 24'sh_051760, 24'sh_0a2c35, 24'sh_144447, 24'sh_27ece1, 24'sh_4b9014, 24'sh_800000 }
