{ 18'sh_00001, 18'sh_00003, 18'sh_00005, 18'sh_0000a, 18'sh_00014, 18'sh_00029, 18'sh_00051, 18'sh_000a3, 18'sh_00146, 18'sh_0028c, 18'sh_00518, 18'sh_00a2f, 18'sh_0145d, 18'sh_028b1, 18'sh_05111, 18'sh_09fb4, 18'sh_12e40, 18'sh_20000 }
